module axi_lite_memory (

);

endmodule


